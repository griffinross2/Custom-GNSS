`ifndef COMMON_GNSS_TYPES_VH
`define COMMON_GNSS_TYPES_VH

// Common types package
package common_gnss_types_pkg;

    typedef logic [4:0] sv_t;
    typedef logic [10:1] l1ca_lfsr_t;
    typedef logic [9:0] chip_t;

endpackage

`endif // COMMON_GNSS_TYPES_VH
